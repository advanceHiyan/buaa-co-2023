`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////
module CMP(GR1,GR2,jump,bpj,op);
input [31:0] GR1,GR2;
input [2:0] op;
output jump,bpj;
assign jump = (GR1 == GR2) ? 1:0;

endmodule
